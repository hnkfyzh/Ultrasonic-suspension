`timescale 1ns/1ps
module speed_setting(
				input clk,	// 50MHz��ʱ��
				input rst_n,	//�͵�ƽ��λ�ź�
				input bps_start,	//���յ����ݺ󣬲�����ʱ�������ź���λ
				output reg clk_bps	// clk_bps�ĸߵ�ƽΪ���ջ��߷�������λ���м������ 
			);

`define BPS_9600
`define CLK_PERIORD	20	//����ʱ������Ϊ20ns(50MHz)
`define BPS_SET		96	//����ͨ�Ų�����Ϊ9600bps(����Ҫ�Ĳ�����ʡȥ��������弴��)

`define BPS_PARA	(10_000_000/`CLK_PERIORD/`BPS_SET)//10_000_000/`CLK_PERIORD/96;		//������Ϊ9600ʱ�ķ�Ƶ����ֵ
`define BPS_PARA_2	(`BPS_PARA/2)//BPS_PARA/2;	//������Ϊ9600ʱ�ķ�Ƶ����ֵ��һ�룬�������ݲ���

reg[15:0] cnt;			//��Ƶ����

//----------------------------------------------------------
reg[2:0] uart_ctrl;	// uart������ѡ��Ĵ���
//----------------------------------------------------------

always @ (posedge clk or negedge rst_n)
	if(!rst_n) cnt <= 16'd0;
	else if((cnt == `BPS_PARA) || !bps_start) cnt <= 16'd0;	//�����ʼ�������
	else cnt <= cnt+1'b1;			//������ʱ�Ӽ�������

always @ (posedge clk or negedge rst_n)
	if(!rst_n) clk_bps <= 1'b0;
	else if(cnt == `BPS_PARA_2) clk_bps <= 1'b1;	// clk_bps_r�ߵ�ƽΪ��������λ���м������,ͬʱҲ��Ϊ�������ݵ����ݸı��
	else clk_bps <= 1'b0;

	
endmodule

